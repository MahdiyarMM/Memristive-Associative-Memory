
.include Models.sp 
.include m.txt
.end